parameter [(2*N_ADD-1):0] COEF_VEC = {2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b11, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b01, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b01, 2'b00, 2'b01, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b01, 2'b00, 2'b00, 2'b00, 2'b11, 2'b00, 2'b00, 2'b00, 2'b00, 2'b11, 2'b00, 2'b00, 2'b00, 2'b11, 2'b00, 2'b00, 2'b11, 2'b00, 2'b00, 2'b00, 2'b00, 2'b01, 2'b00, 2'b00, 2'b00, 2'b11, 2'b00, 2'b00, 2'b01, 2'b00, 2'b00, 2'b11, 2'b00, 2'b00, 2'b00, 2'b11, 2'b00, 2'b01, 2'b00, 2'b01, 2'b00, 2'b11, 2'b00, 2'b00, 2'b00, 2'b00, 2'b01, 2'b00, 2'b00, 2'b11, 2'b00, 2'b00, 2'b00, 2'b11, 2'b00, 2'b00, 2'b00, 2'b01, 2'b00, 2'b00, 2'b00, 2'b11, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b11, 2'b00, 2'b00, 2'b11, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b11, 2'b00, 2'b00, 2'b00, 2'b00, 2'b11, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b01, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b01, 2'b00, 2'b01, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b01, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b11};