* LMV116 - Rev. A
* Created by Bala Ravi; April 16, 2020
* Created with Green-Williams-Lis Op Amp Macro-model Architecture
* Copyright 2020 by Texas Instruments Corporation
******************************************************
* MACRO-MODEL SIMULATED PARAMETERS:
******************************************************
* OPEN-LOOP GAIN AND PHASE VS. FREQUENCY  WITH RL, CL EFFECTS (Aol)
* UNITY GAIN BANDWIDTH (GBW)
* INPUT COMMON-MODE REJECTION RATIO VS. FREQUENCY (CMRR)
* POWER SUPPLY REJECTION RATIO VS. FREQUENCY (PSRR)
* DIFFERENTIAL INPUT IMPEDANCE (Zid)
* COMMON-MODE INPUT IMPEDANCE (Zic)
* OPEN-LOOP OUTPUT IMPEDANCE VS. FREQUENCY (Zo)
* OUTPUT CURRENT THROUGH THE SUPPLY (Iout)
* INPUT VOLTAGE NOISE DENSITY VS. FREQUENCY (en)
* INPUT CURRENT NOISE DENSITY VS. FREQUENCY (in)
* OUTPUT VOLTAGE SWING vs. OUTPUT CURRENT (Vo)
* SHORT-CIRCUIT OUTPUT CURRENT (Isc)
* QUIESCENT CURRENT (Iq)
* SETTLING TIME VS. CAPACITIVE LOAD (ts)
* SLEW RATE (SR)
* SMALL SIGNAL OVERSHOOT VS. CAPACITIVE LOAD
* LARGE SIGNAL RESPONSE
* OVERLOAD RECOVERY TIME (tor)
* INPUT BIAS CURRENT (Ib)
* INPUT OFFSET CURRENT (Ios)
* INPUT OFFSET VOLTAGE (Vos)
* INPUT COMMON-MODE VOLTAGE RANGE (Vcm)
* INPUT OFFSET VOLTAGE VS. INPUT COMMON-MODE VOLTAGE (Vos vs. Vcm)
* INPUT/OUTPUT ESD CELLS (ESDin, ESDout)
******************************************************
.subckt LMV116 IN+ IN- VCC VEE OUT
******************************************************
* MODEL DEFINITIONS:
.model BB_SW VSWITCH(Ron=50 Roff=1e12 Von=700e-3 Voff=0)
.model ESD_SW VSWITCH(Ron=50 Roff=1e12 Von=250e-3 Voff=0)
.model OL_SW VSWITCH(Ron=1e-3 Roff=1e9 Von=900e-3 Voff=800e-3)
.model OR_SW VSWITCH(Ron=10e-3 Roff=1e9 Von=1e-3 Voff=0)
.model R_NOISELESS RES(T_ABS=-273.15)
******************************************************


I_OS        ESDn MID 397N
I_B         23 MID 400N
V_GRp       53 MID 40
V_GRn       54 MID -40
V_ISCp      47 MID 35
V_ISCn      48 MID -32
V_ORn       31 VCLP -80
V11         52 30 0
V_ORp       29 VCLP 80
V12         51 28 0
V4          42 OUT 0
VCM_MIN     75 VEE_B -300M
VCM_MAX     76 VCC_B -1
I_Q         VCC VEE 600U
V_OS        83 23 822.2U
Rsrc        MID 21 R_NOISELESS 1 
G_adjust    21 MID ESDp MID  -148.7M
R48         21 22 R_NOISELESS 100MEG 
C14         22 21 79.58F 
R49         MID 22 R_NOISELESS 44.46K 
SW11        ESDp ESDn ESDp ESDn  S_VSWITCH_1
SW10        ESDn ESDp ESDn ESDp  S_VSWITCH_2
S5          VEE ESDp VEE ESDp  S_VSWITCH_3
S4          VEE ESDn VEE ESDn  S_VSWITCH_4
S2          ESDn VCC ESDn VCC  S_VSWITCH_5
S3          ESDp VCC ESDp VCC  S_VSWITCH_6
C28         24 MID 1P 
R77         25 24 R_NOISELESS 100 
C27         26 MID 1P 
R76         27 26 R_NOISELESS 100 
R75         MID 28 R_NOISELESS 1 
GVCCS8      28 MID 29 MID  -1
R74         30 MID R_NOISELESS 1 
GVCCS7      30 MID 31 MID  -1
R73         32 MID R_NOISELESS 1 
XVCCS_LIM_ZO 33 MID MID 32 VCCS_LIM_ZO_0
Xi_nn       ESDn MID FEMT_0
Xi_np       MID 23 FEMT_0
Xe_n        ESDp 23 VNSE_0
C25         34 MID 3.183F 
R69         MID 34 R_NOISELESS 1MEG 
GVCCS6      34 MID VSENSE MID  -1U
C20         CLAMP MID 125P 
R68         MID CLAMP R_NOISELESS 1MEG 
XVCCS_LIM_2 35 MID MID CLAMP VCCS_LIM_2_0
R44         MID 35 R_NOISELESS 1MEG 
XVCCS_LIM_1 36 37 MID 35 VCCS_LIM_1_0
R72         33 MID R_NOISELESS 2.5 
C26         33 38 63.66F 
R71         33 38 R_NOISELESS 10K 
R70         38 MID R_NOISELESS 1 
GVCCS5      38 MID 39 MID  -1
C23         40 MID 31.83F 
R67         39 40 R_NOISELESS 10K 
R66         39 41 R_NOISELESS 323.3K 
R65         41 MID R_NOISELESS 1 
Rdummy      MID 42 R_NOISELESS 2K 
Rx          42 32 R_NOISELESS 20K 
G_Aol_Zo    41 MID CL_CLAMP 42  -390
R61         MID 43 R_NOISELESS 4.45K 
C16         43 44 795.8F 
R58         44 43 R_NOISELESS 100MEG 
GVCCS2      44 MID VEE_B MID  -471.7M
R57         MID 44 R_NOISELESS 1 
R56         MID 45 R_NOISELESS 10K 
C15         45 46 397.9F 
R55         46 45 R_NOISELESS 100MEG 
GVCCS1      46 MID VCC_B MID  -142.7M
R54         MID 46 R_NOISELESS 1 
XIQPos      VIMON MID MID VCC VCCS_LIMIT_IQ_0
XIQNeg      MID VIMON VEE MID VCCS_LIMIT_IQ_0
C_DIFF      ESDp ESDn 4P 
XCL_AMP     47 48 VIMON MID 49 50 CLAMP_AMP_LO_0
SOR_SWp     CLAMP 51 CLAMP 51  S_VSWITCH_7
SOR_SWn     52 CLAMP 52 CLAMP  S_VSWITCH_8
XGR_AMP     53 54 55 MID 56 57 CLAMP_AMP_HI_0
R39         53 MID R_NOISELESS 1T 
R37         54 MID R_NOISELESS 1T 
R42         VSENSE 55 R_NOISELESS 1M 
C19         55 MID 1F 
R38         56 MID R_NOISELESS 1 
R36         MID 57 R_NOISELESS 1 
R40         56 58 R_NOISELESS 1M 
R41         57 59 R_NOISELESS 1M 
C17         58 MID 1F 
C18         MID 59 1F 
XGR_SRC     58 59 CLAMP MID VCCS_LIM_GR_0
R21         49 MID R_NOISELESS 1 
R20         MID 50 R_NOISELESS 1 
R29         49 60 R_NOISELESS 1M 
R30         50 61 R_NOISELESS 1M 
C9          60 MID 1F 
C8          MID 61 1F 
XCL_SRC     60 61 CL_CLAMP MID VCCS_LIM_4_0
R22         47 MID R_NOISELESS 1T 
R19         MID 48 R_NOISELESS 1T 
XCLAWp      VIMON MID 62 VCC_B VCCS_LIM_CLAW+_0
XCLAWn      MID VIMON VEE_B 63 VCCS_LIM_CLAW-_0
R12         62 VCC_B R_NOISELESS 1K 
R16         62 64 R_NOISELESS 1M 
R13         VEE_B 63 R_NOISELESS 1K 
R17         65 63 R_NOISELESS 1M 
C6          65 MID 1F 
C5          MID 64 1F 
G2          VCC_CLP MID 64 MID  -1M
R15         VCC_CLP MID R_NOISELESS 1K 
G3          VEE_CLP MID 65 MID  -1M
R14         MID VEE_CLP R_NOISELESS 1K 
XCLAW_AMP   VCC_CLP VEE_CLP VOUT_S MID 66 67 CLAMP_AMP_LO_0
R26         VCC_CLP MID R_NOISELESS 1T 
R23         VEE_CLP MID R_NOISELESS 1T 
R25         66 MID R_NOISELESS 1 
R24         MID 67 R_NOISELESS 1 
R27         66 68 R_NOISELESS 1M 
R28         67 69 R_NOISELESS 1M 
C11         68 MID 1F 
C10         MID 69 1F 
XCLAW_SRC   68 69 CLAW_CLAMP MID VCCS_LIM_3_0
H2          27 MID V11 -1
H3          25 MID V12 1
C12         SW_OL MID 100P 
R32         70 SW_OL R_NOISELESS 100 
R31         70 MID R_NOISELESS 1 
XOL_SENSE   MID 70 26 24 OL_SENSE_0
S1          41 39 SW_OL MID  S_VSWITCH_9
H1          71 MID V4 1K
S7          VEE OUT VEE OUT  S_VSWITCH_10
S6          OUT VCC OUT VCC  S_VSWITCH_11
R11         MID 72 R_NOISELESS 1T 
R18         72 VOUT_S R_NOISELESS 100 
C7          VOUT_S MID 1N 
E5          72 MID OUT MID  1
C13         VIMON MID 1N 
R33         71 VIMON R_NOISELESS 100 
R10         MID 71 R_NOISELESS 1T 
R47         73 VCLP R_NOISELESS 100 
C24         VCLP MID 100P 
E4          73 MID CL_CLAMP MID  1
R46         MID CL_CLAMP R_NOISELESS 1K 
G9          CL_CLAMP MID CLAW_CLAMP MID  -1M
R45         MID CLAW_CLAMP R_NOISELESS 1K 
G8          CLAW_CLAMP MID 34 MID  -1M
R43         MID VSENSE R_NOISELESS 1K 
G15         VSENSE MID CLAMP MID  -1M
C4          36 MID 1F 
R9          36 74 R_NOISELESS 1M 
R7          MID 75 R_NOISELESS 1T 
R6          76 MID R_NOISELESS 1T 
R8          MID 74 R_NOISELESS 1 
XVCM_CLAMP  77 MID 74 MID 76 75 VCCS_EXT_LIM_0
E1          MID 0 78 0  1
R89         VEE_B 0 R_NOISELESS 1 
R5          79 VEE_B R_NOISELESS 1M 
C3          79 0 1F 
R60         78 79 R_NOISELESS 1MEG 
C1          78 0 1 
R3          78 0 R_NOISELESS 1T 
R59         80 78 R_NOISELESS 1MEG 
C2          80 0 1F 
R4          VCC_B 80 R_NOISELESS 1M 
R88         VCC_B 0 R_NOISELESS 1 
G17         VEE_B 0 VEE 0  -1
G16         VCC_B 0 VCC 0  -1
R_PSR       81 77 R_NOISELESS 1K 
G_PSR       77 81 45 43  -1M
R2          37 ESDn R_NOISELESS 1M 
R1          81 82 R_NOISELESS 1M 
R_CMR       83 82 R_NOISELESS 1K 
G_CMR       82 83 22 MID  -1M
C_CMn       ESDn MID 2P 
C_CMp       MID ESDp 2P 
R53         ESDn MID R_NOISELESS 1T 
R52         MID ESDp R_NOISELESS 1T 
R35         IN- ESDn R_NOISELESS 10M 
R34         IN+ ESDp R_NOISELESS 10M 

.MODEL S_VSWITCH_1 VSWITCH (RON=50 ROFF=1T VON=700M VOFF=0)
.MODEL S_VSWITCH_2 VSWITCH (RON=50 ROFF=1T VON=700M VOFF=0)
.MODEL S_VSWITCH_3 VSWITCH (RON=50 ROFF=1T VON=500M VOFF=100M)
.MODEL S_VSWITCH_4 VSWITCH (RON=50 ROFF=1T VON=500M VOFF=100M)
.MODEL S_VSWITCH_5 VSWITCH (RON=50 ROFF=1T VON=500M VOFF=100M)
.MODEL S_VSWITCH_6 VSWITCH (RON=50 ROFF=1T VON=500M VOFF=100M)
.MODEL S_VSWITCH_7 VSWITCH (RON=10M ROFF=1T VON=10M VOFF=0)
.MODEL S_VSWITCH_8 VSWITCH (RON=10M ROFF=1T VON=10M VOFF=0)
.MODEL S_VSWITCH_9 VSWITCH (RON=1M ROFF=1T VON=500M VOFF=100M)
.MODEL S_VSWITCH_10 VSWITCH (RON=50 ROFF=1T VON=500M VOFF=100M)
.MODEL S_VSWITCH_11 VSWITCH (RON=50 ROFF=1T VON=500M VOFF=100M)

.ENDS LMV116
*
.SUBCKT VCCS_LIM_ZO_0  VC+ VC- IOUT+ IOUT-
.PARAM GAIN = 4E3
.PARAM IPOS = 1E6
.PARAM INEG = -1E6
G1 IOUT+ IOUT- VALUE={LIMIT(GAIN*V(VC+,VC-),INEG,IPOS)}
.ENDS
*


.SUBCKT FEMT_0  1 2
.PARAM FLWF=10
.PARAM NLFF=4500
.PARAM NVRF=750
.PARAM GLFF={PWR(FLWF,0.25)*NLFF/1164}
.PARAM RNVF={1.184*PWR(NVRF,2)}
.MODEL DVNF D KF={PWR(FLWF,0.5)/1E11} IS=1.0E-16
I1 0 7 10E-3
I2 0 8 10E-3
D1 7 0 DVNF
D2 8 0 DVNF
E1 3 6 7 8 {GLFF}
R1 3 0 1E9
R2 3 0 1E9
R3 3 6 1E9
E2 6 4 5 0 10
R4 5 0 {RNVF}
R5 5 0 {RNVF}
R6 3 4 1E9
R7 4 0 1E9
G1 1 2 3 4 1E-6
.ENDS
*


.SUBCKT VNSE_0  1 2
.PARAM FLW=10
.PARAM NLF=450
.PARAM NVR=35
.PARAM GLF={PWR(FLW,0.25)*NLF/1164}
.PARAM RNV={1.184*PWR(NVR,2)}
.MODEL DVN D KF={PWR(FLW,0.5)/1E11} IS=1.0E-16
I1 0 7 10E-3
I2 0 8 10E-3
D1 7 0 DVN
D2 8 0 DVN
E1 3 6 7 8 {GLF}
R1 3 0 1E9
R2 3 0 1E9
R3 3 6 1E9
E2 6 4 5 0 10
R4 5 0 {RNV}
R5 5 0 {RNV}
R6 3 4 1E9
R7 4 0 1E9
E3 1 2 3 4 1
.ENDS
*


.SUBCKT VCCS_LIM_2_0  VC+ VC- IOUT+ IOUT-
.PARAM GAIN = 3.32E-4
.PARAM IPOS = 0.005
.PARAM INEG = -0.005
G1 IOUT+ IOUT- VALUE={LIMIT(GAIN*V(VC+,VC-),INEG,IPOS)}
.ENDS
*



.SUBCKT VCCS_LIM_1_0  VC+ VC- IOUT+ IOUT-
.PARAM GAIN = 1E-4
.PARAM IPOS = .5
.PARAM INEG = -.5
G1 IOUT+ IOUT- VALUE={LIMIT(GAIN*V(VC+,VC-),INEG,IPOS)}
.ENDS
*


.SUBCKT VCCS_LIMIT_IQ_0  VC+ VC- IOUT+ IOUT-
.PARAM GAIN = 1E-3
G1 IOUT- IOUT+ VALUE={IF( (V(VC+,VC-)<=0),0,GAIN*V(VC+,VC-) )}
.ENDS
*


.SUBCKT CLAMP_AMP_LO_0  VC+ VC- VIN COM VO+ VO-
.PARAM G=1
GVO+ COM VO+ VALUE = {IF(V(VIN,COM)>V(VC+,COM),((V(VIN,COM)-V(VC+,COM))*G),0)}
GVO- COM VO- VALUE = {IF(V(VIN,COM)<V(VC-,COM),((V(VC-,COM)-V(VIN,COM))*G),0)}
.ENDS
*


.SUBCKT CLAMP_AMP_HI_0  VC+ VC- VIN COM VO+ VO-
.PARAM G=10
GVO+ COM VO+ VALUE = {IF(V(VIN,COM)>V(VC+,COM),((V(VIN,COM)-V(VC+,COM))*G),0)}
GVO- COM VO- VALUE = {IF(V(VIN,COM)<V(VC-,COM),((V(VC-,COM)-V(VIN,COM))*G),0)}
.ENDS
*


.SUBCKT VCCS_LIM_GR_0  VC+ VC- IOUT+ IOUT-
.PARAM GAIN = 1
.PARAM IPOS = 11
.PARAM INEG = -11
G1 IOUT+ IOUT- VALUE={LIMIT(GAIN*V(VC+,VC-),INEG,IPOS)}
.ENDS
*


.SUBCKT VCCS_LIM_4_0  VC+ VC- IOUT+ IOUT-
.PARAM GAIN = 1
.PARAM IPOS = 550E-3
.PARAM INEG = -550E-3
G1 IOUT+ IOUT- VALUE={LIMIT(GAIN*V(VC+,VC-),INEG,IPOS)}
.ENDS
*


.SUBCKT VCCS_LIM_CLAW+_0  VC+ VC- IOUT+ IOUT-
G1 IOUT+ IOUT- TABLE {ABS(V(VC+,VC-))} =
+(0, 1E-5)
+(10.52, 1.2E-4)
+(20.45, 2.2E-4)
+(28.244, 3.46E-4)
+(34.42, 8.23E-4)
+(39.74, 1.6E-3)
+(43.8, 2.4E-3)
.ENDS
*


.SUBCKT VCCS_LIM_CLAW-_0  VC+ VC- IOUT+ IOUT-
G1 IOUT+ IOUT- TABLE {ABS(V(VC+,VC-))} =
+(0, 5E-5)
+(25, 4E-4)
+(29, 5.67E-4)
+(32.2, 8.2E-4)
+(38.11, 1.68E-3)
+(40.25, 2.09E-3)
+(42.23, 2.5E-3)
.ENDS
*


.SUBCKT VCCS_LIM_3_0  VC+ VC- IOUT+ IOUT-
.PARAM GAIN = 1
.PARAM IPOS = 530E-3
.PARAM INEG = -530E-3
G1 IOUT+ IOUT- VALUE={LIMIT(GAIN*V(VC+,VC-),INEG,IPOS)}
.ENDS
*


.SUBCKT OL_SENSE_0  COM SW+ OLN  OLP
GSW+ COM SW+ VALUE = {IF((V(OLN,COM)>10E-3 | V(OLP,COM)>10E-3),1,0)}
.ENDS
*


.SUBCKT VCCS_EXT_LIM_0  VIN+ VIN- IOUT- IOUT+ VP+ VP-
.PARAM GAIN = 1
G1 IOUT+ IOUT- VALUE={LIMIT(GAIN*V(VIN+,VIN-),V(VP-,VIN-), V(VP+,VIN-))}
.ENDS
*


